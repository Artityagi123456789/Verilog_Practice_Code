//XNOR Gate Design File
module XNOR(input a,b, output out);
  xnor G(out,a,b);
endmodule


